typedef enum logic [2:0] {
  // Will be added when implementing the operations
} alu_operation_e;
